module encoder 
#(parameter bits = 8,
parameter stages = 10)(
    input clk,
    input rst,
    input [9:0] data,
    output reg [7:0] encoded_data
);



endmodule
